module (
    input SDRAM_EN,
    input CLK,
    input RST_L,
    input [3:0] SDRAM_CYCLE,
    input [3:0] STATE_CNTR,
    output [11:0] SDRAM_MODE_REG,
    output [1:0] SDRAM_CMND,
    output CMND_CYCE_REQ,
    output SDRAM_SETUP
);

//Add logic here





endmodule
