module (
    input CLK,
    input RST_L,
    input SDRAM_SETUP,
    input [3:0] SDRAM_CYCLE,
    output RFRSH_REQ
);

//Add logic here





endmodule
