module (
    input CLK,
    input SDRAM_CS_L,
    input CMND_CYCL_REQ,
    input RFRSH_REQ,
    input RST_L,
    output SDRAM_CYCLE,
    output [3:0] STATE_CNTR,
);

//Add logic here





endmodule
